/* Verilog model created from schematic DSPmaster.sch -- Jan 15, 2018 14:27 */

module DSPmaster;




endmodule // DSPmaster
